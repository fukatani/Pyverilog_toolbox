module TOP(CLK, RST);
  input CLK,RST;
  wire wire1;

  assign wire1 = wire1;

endmodule

